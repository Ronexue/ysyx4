
module mytest;
initial begin $display("hello world"); end
endmodule
